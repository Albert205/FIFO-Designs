// Code your design here
`include "fifo_ctrl.sv"
`include "fifo_top.sv"
`include "register_file.sv"
`include "interface.sv"